module vga_clock_gen(
	
);