module custom_multiply (
	
	// Inputs required for multicycle custom instructions

	input [31:0] dataa,
	input [31:0] datab,

	// Outputs
	output [31:0] result

);

always @(posedge clk or posedge reset) begin
    
end
